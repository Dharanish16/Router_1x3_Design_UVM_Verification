
module router_sync(clock,resetn,data_in,detect_add,full_0,full_1,full_2,empty_0,
                   empty_1,empty_2,write_enb_reg,read_enb_0,read_enb_1,
						 read_enb_2,vld_out_0,vld_out_1,vld_out_2,fifo_full,
						 soft_reset_0,soft_reset_1,soft_reset_2,write_enb);
        input [1:0]data_in;
		  input clock,resetn,detect_add,full_0,full_1,full_2,empty_0,empty_1,empty_2,write_enb_reg,read_enb_0,read_enb_1,read_enb_2;
		  output vld_out_0,vld_out_1,vld_out_2;
		  output reg soft_reset_0,soft_reset_1,soft_reset_2;
		  output reg[2:0]write_enb;
		  output reg fifo_full;
		  reg [1:0]temp;
		  reg [4:0]count0,count1,count2;
		  
		  
		  //RTL schematic for capturing address
		  always@(posedge clock)
		      begin
				   if(!resetn)
					   temp <= 0;
				   else if(detect_add)
					   temp <= data_in;
					else 
					   temp <= temp;
			   end
		  
		  //fifo_full logic using case statement
		  always@(*)
		      begin
				   case(temp)
					    2'b00 : fifo_full = full_0;
						 2'b01 : fifo_full = full_1;
						 2'b10 : fifo_full = full_2;
						 default : fifo_full = 0;
					endcase
			   end
				
			//write enable logic
			always@(*)
			    begin
				    if(write_enb_reg)
					     begin
						     case(temp)
							      2'b00  :  write_enb = 3'b001;
									2'b01  :  write_enb = 3'b010;
									2'b10  :  write_enb = 3'b100;
									default : write_enb = 3'b000;
							  endcase
						  end
					 else
					    write_enb = 3'b000;
				end
		  
		   //Direct assignment for valid out signals
			assign vld_out_0 = ~empty_0;
			assign vld_out_1 = ~empty_1;
			assign vld_out_2 = ~empty_2;
			
			//Logic for soft_reset_0
			always@(posedge clock)
			    begin
				     if(!resetn)
					        count0 <= 5'b0;
					  else if(vld_out_0)
					     begin
						     if(!read_enb_0)
									begin
										if(count0 == 5'd29)
												begin
													soft_reset_0 <= 1'b1;
													count0 <= 5'b0;
												end
										else
												begin
													count0 <= count0 + 5'b1;
													soft_reset_0 <= 1'b0;
												end
									end
							   else
									count0 <= 5'b0;
						  end
					  else
					    count0 <= 5'b0;
				  end
				  
			//Logic for soft_reset_1
			always@(posedge clock)
			    begin
				     if(!resetn)
					        count1 <= 5'b0;
					  else if(vld_out_1)
					     begin
						     if(!read_enb_1)
									begin
										if(count1 == 5'd29)
												begin
													soft_reset_1 <= 1'b1;
													count1 <= 5'b0;
												end
										else
												begin
													count1 <= count1 + 5'b1;
													soft_reset_1 <= 1'b0;
												end
									end
							   else
									count1 <= 5'b0;
						  end
					  else
					    count1 <= 5'b0;
				  end
		    
			//Logic for soft_reset_2
			 always@(posedge clock)
			    begin
				     if(!resetn)
					        count2 <= 5'b0;
					  else if(vld_out_2)
					     begin
						     if(!read_enb_2)
									begin
										if(count2 == 5'd29)
												begin
													soft_reset_2 <= 1'b1;
													count2 <= 5'b0;
												end
										else
												begin
													count2 <= count2 + 5'b1;
													soft_reset_2 <= 1'b0;
												end
									end
							   else
									count2 <= 5'b0;
						  end
					  else
					    count2 <= 5'b0;
				  end
endmodule

							  
			
			
						 